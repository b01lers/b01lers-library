`timescale 1 ns/10 ps  // time-unit = 1 ns, precision = 10 ps

module test;
  reg ENABLE = 0;
  reg RESET = 0;
  reg [127:0] PLAINTEXT = 0;

  initial begin
     # 100 RESET = 1;
     # 100 ENABLE = 0;


     # 200 RESET = 0;
     # 200 ENABLE = 1;

     # 3000 $stop;
  end


    reg CLK = 0;
    initial CLK = 0; 
  always #10 CLK = ~CLK; 

  wire [127:0] CIPHERTEXT;
  wire  DONE;

  AES128 aes128_inst (
    .CLK (CLK),
    .RESET (RESET),
    .ENABLE (ENABLE),
    .DONE (DONE),
    .PLAINTEXT_0 (PLAINTEXT[0]),
    .PLAINTEXT_1 (PLAINTEXT[1]),
    .PLAINTEXT_2 (PLAINTEXT[2]),
    .PLAINTEXT_3 (PLAINTEXT[3]),
    .PLAINTEXT_4 (PLAINTEXT[4]),
    .PLAINTEXT_5 (PLAINTEXT[5]),
    .PLAINTEXT_6 (PLAINTEXT[6]),
    .PLAINTEXT_7 (PLAINTEXT[7]),
    .PLAINTEXT_8 (PLAINTEXT[8]),
    .PLAINTEXT_9 (PLAINTEXT[9]),
    .PLAINTEXT_10 (PLAINTEXT[10]),
    .PLAINTEXT_11 (PLAINTEXT[11]),
    .PLAINTEXT_12 (PLAINTEXT[12]),
    .PLAINTEXT_13 (PLAINTEXT[13]),
    .PLAINTEXT_14 (PLAINTEXT[14]),
    .PLAINTEXT_15 (PLAINTEXT[15]),
    .PLAINTEXT_16 (PLAINTEXT[16]),
    .PLAINTEXT_17 (PLAINTEXT[17]),
    .PLAINTEXT_18 (PLAINTEXT[18]),
    .PLAINTEXT_19 (PLAINTEXT[19]),
    .PLAINTEXT_20 (PLAINTEXT[20]),
    .PLAINTEXT_21 (PLAINTEXT[21]),
    .PLAINTEXT_22 (PLAINTEXT[22]),
    .PLAINTEXT_23 (PLAINTEXT[23]),
    .PLAINTEXT_24 (PLAINTEXT[24]),
    .PLAINTEXT_25 (PLAINTEXT[25]),
    .PLAINTEXT_26 (PLAINTEXT[26]),
    .PLAINTEXT_27 (PLAINTEXT[27]),
    .PLAINTEXT_28 (PLAINTEXT[28]),
    .PLAINTEXT_29 (PLAINTEXT[29]),
    .PLAINTEXT_30 (PLAINTEXT[30]),
    .PLAINTEXT_31 (PLAINTEXT[31]),
    .PLAINTEXT_32 (PLAINTEXT[32]),
    .PLAINTEXT_33 (PLAINTEXT[33]),
    .PLAINTEXT_34 (PLAINTEXT[34]),
    .PLAINTEXT_35 (PLAINTEXT[35]),
    .PLAINTEXT_36 (PLAINTEXT[36]),
    .PLAINTEXT_37 (PLAINTEXT[37]),
    .PLAINTEXT_38 (PLAINTEXT[38]),
    .PLAINTEXT_39 (PLAINTEXT[39]),
    .PLAINTEXT_40 (PLAINTEXT[40]),
    .PLAINTEXT_41 (PLAINTEXT[41]),
    .PLAINTEXT_42 (PLAINTEXT[42]),
    .PLAINTEXT_43 (PLAINTEXT[43]),
    .PLAINTEXT_44 (PLAINTEXT[44]),
    .PLAINTEXT_45 (PLAINTEXT[45]),
    .PLAINTEXT_46 (PLAINTEXT[46]),
    .PLAINTEXT_47 (PLAINTEXT[47]),
    .PLAINTEXT_48 (PLAINTEXT[48]),
    .PLAINTEXT_49 (PLAINTEXT[49]),
    .PLAINTEXT_50 (PLAINTEXT[50]),
    .PLAINTEXT_51 (PLAINTEXT[51]),
    .PLAINTEXT_52 (PLAINTEXT[52]),
    .PLAINTEXT_53 (PLAINTEXT[53]),
    .PLAINTEXT_54 (PLAINTEXT[54]),
    .PLAINTEXT_55 (PLAINTEXT[55]),
    .PLAINTEXT_56 (PLAINTEXT[56]),
    .PLAINTEXT_57 (PLAINTEXT[57]),
    .PLAINTEXT_58 (PLAINTEXT[58]),
    .PLAINTEXT_59 (PLAINTEXT[59]),
    .PLAINTEXT_60 (PLAINTEXT[60]),
    .PLAINTEXT_61 (PLAINTEXT[61]),
    .PLAINTEXT_62 (PLAINTEXT[62]),
    .PLAINTEXT_63 (PLAINTEXT[63]),
    .PLAINTEXT_64 (PLAINTEXT[64]),
    .PLAINTEXT_65 (PLAINTEXT[65]),
    .PLAINTEXT_66 (PLAINTEXT[66]),
    .PLAINTEXT_67 (PLAINTEXT[67]),
    .PLAINTEXT_68 (PLAINTEXT[68]),
    .PLAINTEXT_69 (PLAINTEXT[69]),
    .PLAINTEXT_70 (PLAINTEXT[70]),
    .PLAINTEXT_71 (PLAINTEXT[71]),
    .PLAINTEXT_72 (PLAINTEXT[72]),
    .PLAINTEXT_73 (PLAINTEXT[73]),
    .PLAINTEXT_74 (PLAINTEXT[74]),
    .PLAINTEXT_75 (PLAINTEXT[75]),
    .PLAINTEXT_76 (PLAINTEXT[76]),
    .PLAINTEXT_77 (PLAINTEXT[77]),
    .PLAINTEXT_78 (PLAINTEXT[78]),
    .PLAINTEXT_79 (PLAINTEXT[79]),
    .PLAINTEXT_80 (PLAINTEXT[80]),
    .PLAINTEXT_81 (PLAINTEXT[81]),
    .PLAINTEXT_82 (PLAINTEXT[82]),
    .PLAINTEXT_83 (PLAINTEXT[83]),
    .PLAINTEXT_84 (PLAINTEXT[84]),
    .PLAINTEXT_85 (PLAINTEXT[85]),
    .PLAINTEXT_86 (PLAINTEXT[86]),
    .PLAINTEXT_87 (PLAINTEXT[87]),
    .PLAINTEXT_88 (PLAINTEXT[88]),
    .PLAINTEXT_89 (PLAINTEXT[89]),
    .PLAINTEXT_90 (PLAINTEXT[90]),
    .PLAINTEXT_91 (PLAINTEXT[91]),
    .PLAINTEXT_92 (PLAINTEXT[92]),
    .PLAINTEXT_93 (PLAINTEXT[93]),
    .PLAINTEXT_94 (PLAINTEXT[94]),
    .PLAINTEXT_95 (PLAINTEXT[95]),
    .PLAINTEXT_96 (PLAINTEXT[96]),
    .PLAINTEXT_97 (PLAINTEXT[97]),
    .PLAINTEXT_98 (PLAINTEXT[98]),
    .PLAINTEXT_99 (PLAINTEXT[99]),
    .PLAINTEXT_100 (PLAINTEXT[100]),
    .PLAINTEXT_101 (PLAINTEXT[101]),
    .PLAINTEXT_102 (PLAINTEXT[102]),
    .PLAINTEXT_103 (PLAINTEXT[103]),
    .PLAINTEXT_104 (PLAINTEXT[104]),
    .PLAINTEXT_105 (PLAINTEXT[105]),
    .PLAINTEXT_106 (PLAINTEXT[106]),
    .PLAINTEXT_107 (PLAINTEXT[107]),
    .PLAINTEXT_108 (PLAINTEXT[108]),
    .PLAINTEXT_109 (PLAINTEXT[109]),
    .PLAINTEXT_110 (PLAINTEXT[110]),
    .PLAINTEXT_111 (PLAINTEXT[111]),
    .PLAINTEXT_112 (PLAINTEXT[112]),
    .PLAINTEXT_113 (PLAINTEXT[113]),
    .PLAINTEXT_114 (PLAINTEXT[114]),
    .PLAINTEXT_115 (PLAINTEXT[115]),
    .PLAINTEXT_116 (PLAINTEXT[116]),
    .PLAINTEXT_117 (PLAINTEXT[117]),
    .PLAINTEXT_118 (PLAINTEXT[118]),
    .PLAINTEXT_119 (PLAINTEXT[119]),
    .PLAINTEXT_120 (PLAINTEXT[120]),
    .PLAINTEXT_121 (PLAINTEXT[121]),
    .PLAINTEXT_122 (PLAINTEXT[122]),
    .PLAINTEXT_123 (PLAINTEXT[123]),
    .PLAINTEXT_124 (PLAINTEXT[124]),
    .PLAINTEXT_125 (PLAINTEXT[125]),
    .PLAINTEXT_126 (PLAINTEXT[126]),
    .PLAINTEXT_127 (PLAINTEXT[127]),
    .CIPHERTEXT_0 (CIPHERTEXT[0]),
    .CIPHERTEXT_1 (CIPHERTEXT[1]),
    .CIPHERTEXT_2 (CIPHERTEXT[2]),
    .CIPHERTEXT_3 (CIPHERTEXT[3]),
    .CIPHERTEXT_4 (CIPHERTEXT[4]),
    .CIPHERTEXT_5 (CIPHERTEXT[5]),
    .CIPHERTEXT_6 (CIPHERTEXT[6]),
    .CIPHERTEXT_7 (CIPHERTEXT[7]),
    .CIPHERTEXT_8 (CIPHERTEXT[8]),
    .CIPHERTEXT_9 (CIPHERTEXT[9]),
    .CIPHERTEXT_10 (CIPHERTEXT[10]),
    .CIPHERTEXT_11 (CIPHERTEXT[11]),
    .CIPHERTEXT_12 (CIPHERTEXT[12]),
    .CIPHERTEXT_13 (CIPHERTEXT[13]),
    .CIPHERTEXT_14 (CIPHERTEXT[14]),
    .CIPHERTEXT_15 (CIPHERTEXT[15]),
    .CIPHERTEXT_16 (CIPHERTEXT[16]),
    .CIPHERTEXT_17 (CIPHERTEXT[17]),
    .CIPHERTEXT_18 (CIPHERTEXT[18]),
    .CIPHERTEXT_19 (CIPHERTEXT[19]),
    .CIPHERTEXT_20 (CIPHERTEXT[20]),
    .CIPHERTEXT_21 (CIPHERTEXT[21]),
    .CIPHERTEXT_22 (CIPHERTEXT[22]),
    .CIPHERTEXT_23 (CIPHERTEXT[23]),
    .CIPHERTEXT_24 (CIPHERTEXT[24]),
    .CIPHERTEXT_25 (CIPHERTEXT[25]),
    .CIPHERTEXT_26 (CIPHERTEXT[26]),
    .CIPHERTEXT_27 (CIPHERTEXT[27]),
    .CIPHERTEXT_28 (CIPHERTEXT[28]),
    .CIPHERTEXT_29 (CIPHERTEXT[29]),
    .CIPHERTEXT_30 (CIPHERTEXT[30]),
    .CIPHERTEXT_31 (CIPHERTEXT[31]),
    .CIPHERTEXT_32 (CIPHERTEXT[32]),
    .CIPHERTEXT_33 (CIPHERTEXT[33]),
    .CIPHERTEXT_34 (CIPHERTEXT[34]),
    .CIPHERTEXT_35 (CIPHERTEXT[35]),
    .CIPHERTEXT_36 (CIPHERTEXT[36]),
    .CIPHERTEXT_37 (CIPHERTEXT[37]),
    .CIPHERTEXT_38 (CIPHERTEXT[38]),
    .CIPHERTEXT_39 (CIPHERTEXT[39]),
    .CIPHERTEXT_40 (CIPHERTEXT[40]),
    .CIPHERTEXT_41 (CIPHERTEXT[41]),
    .CIPHERTEXT_42 (CIPHERTEXT[42]),
    .CIPHERTEXT_43 (CIPHERTEXT[43]),
    .CIPHERTEXT_44 (CIPHERTEXT[44]),
    .CIPHERTEXT_45 (CIPHERTEXT[45]),
    .CIPHERTEXT_46 (CIPHERTEXT[46]),
    .CIPHERTEXT_47 (CIPHERTEXT[47]),
    .CIPHERTEXT_48 (CIPHERTEXT[48]),
    .CIPHERTEXT_49 (CIPHERTEXT[49]),
    .CIPHERTEXT_50 (CIPHERTEXT[50]),
    .CIPHERTEXT_51 (CIPHERTEXT[51]),
    .CIPHERTEXT_52 (CIPHERTEXT[52]),
    .CIPHERTEXT_53 (CIPHERTEXT[53]),
    .CIPHERTEXT_54 (CIPHERTEXT[54]),
    .CIPHERTEXT_55 (CIPHERTEXT[55]),
    .CIPHERTEXT_56 (CIPHERTEXT[56]),
    .CIPHERTEXT_57 (CIPHERTEXT[57]),
    .CIPHERTEXT_58 (CIPHERTEXT[58]),
    .CIPHERTEXT_59 (CIPHERTEXT[59]),
    .CIPHERTEXT_60 (CIPHERTEXT[60]),
    .CIPHERTEXT_61 (CIPHERTEXT[61]),
    .CIPHERTEXT_62 (CIPHERTEXT[62]),
    .CIPHERTEXT_63 (CIPHERTEXT[63]),
    .CIPHERTEXT_64 (CIPHERTEXT[64]),
    .CIPHERTEXT_65 (CIPHERTEXT[65]),
    .CIPHERTEXT_66 (CIPHERTEXT[66]),
    .CIPHERTEXT_67 (CIPHERTEXT[67]),
    .CIPHERTEXT_68 (CIPHERTEXT[68]),
    .CIPHERTEXT_69 (CIPHERTEXT[69]),
    .CIPHERTEXT_70 (CIPHERTEXT[70]),
    .CIPHERTEXT_71 (CIPHERTEXT[71]),
    .CIPHERTEXT_72 (CIPHERTEXT[72]),
    .CIPHERTEXT_73 (CIPHERTEXT[73]),
    .CIPHERTEXT_74 (CIPHERTEXT[74]),
    .CIPHERTEXT_75 (CIPHERTEXT[75]),
    .CIPHERTEXT_76 (CIPHERTEXT[76]),
    .CIPHERTEXT_77 (CIPHERTEXT[77]),
    .CIPHERTEXT_78 (CIPHERTEXT[78]),
    .CIPHERTEXT_79 (CIPHERTEXT[79]),
    .CIPHERTEXT_80 (CIPHERTEXT[80]),
    .CIPHERTEXT_81 (CIPHERTEXT[81]),
    .CIPHERTEXT_82 (CIPHERTEXT[82]),
    .CIPHERTEXT_83 (CIPHERTEXT[83]),
    .CIPHERTEXT_84 (CIPHERTEXT[84]),
    .CIPHERTEXT_85 (CIPHERTEXT[85]),
    .CIPHERTEXT_86 (CIPHERTEXT[86]),
    .CIPHERTEXT_87 (CIPHERTEXT[87]),
    .CIPHERTEXT_88 (CIPHERTEXT[88]),
    .CIPHERTEXT_89 (CIPHERTEXT[89]),
    .CIPHERTEXT_90 (CIPHERTEXT[90]),
    .CIPHERTEXT_91 (CIPHERTEXT[91]),
    .CIPHERTEXT_92 (CIPHERTEXT[92]),
    .CIPHERTEXT_93 (CIPHERTEXT[93]),
    .CIPHERTEXT_94 (CIPHERTEXT[94]),
    .CIPHERTEXT_95 (CIPHERTEXT[95]),
    .CIPHERTEXT_96 (CIPHERTEXT[96]),
    .CIPHERTEXT_97 (CIPHERTEXT[97]),
    .CIPHERTEXT_98 (CIPHERTEXT[98]),
    .CIPHERTEXT_99 (CIPHERTEXT[99]),
    .CIPHERTEXT_100 (CIPHERTEXT[100]),
    .CIPHERTEXT_101 (CIPHERTEXT[101]),
    .CIPHERTEXT_102 (CIPHERTEXT[102]),
    .CIPHERTEXT_103 (CIPHERTEXT[103]),
    .CIPHERTEXT_104 (CIPHERTEXT[104]),
    .CIPHERTEXT_105 (CIPHERTEXT[105]),
    .CIPHERTEXT_106 (CIPHERTEXT[106]),
    .CIPHERTEXT_107 (CIPHERTEXT[107]),
    .CIPHERTEXT_108 (CIPHERTEXT[108]),
    .CIPHERTEXT_109 (CIPHERTEXT[109]),
    .CIPHERTEXT_110 (CIPHERTEXT[110]),
    .CIPHERTEXT_111 (CIPHERTEXT[111]),
    .CIPHERTEXT_112 (CIPHERTEXT[112]),
    .CIPHERTEXT_113 (CIPHERTEXT[113]),
    .CIPHERTEXT_114 (CIPHERTEXT[114]),
    .CIPHERTEXT_115 (CIPHERTEXT[115]),
    .CIPHERTEXT_116 (CIPHERTEXT[116]),
    .CIPHERTEXT_117 (CIPHERTEXT[117]),
    .CIPHERTEXT_118 (CIPHERTEXT[118]),
    .CIPHERTEXT_119 (CIPHERTEXT[119]),
    .CIPHERTEXT_120 (CIPHERTEXT[120]),
    .CIPHERTEXT_121 (CIPHERTEXT[121]),
    .CIPHERTEXT_122 (CIPHERTEXT[122]),
    .CIPHERTEXT_123 (CIPHERTEXT[123]),
    .CIPHERTEXT_124 (CIPHERTEXT[124]),
    .CIPHERTEXT_125 (CIPHERTEXT[125]),
    .CIPHERTEXT_126 (CIPHERTEXT[126]),
    .CIPHERTEXT_127 (CIPHERTEXT[127]));

  initial
     $monitor("At time %t, value = %h (%0d)",
              $time, CIPHERTEXT, CIPHERTEXT);
endmodule // test

